`include "R2/alu.sv"
`include "R2/mux.sv"
`include "R2/regFile.sv"
`include "R3/cu.sv"
`include "R3/ext32.sv"
`include "R3/rom.sv"

module top(
    input wire clk,
    input wire rst,
    output wire a0
);



endmodule
