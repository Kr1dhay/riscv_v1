module 2_ALU(
    input logic 
);