module alu_2 (
    input logic [31:0] aluOp1,
    input logic [31:0] aluOp2,
    input logic [2:0] aluCTR,
    output logic [31:0] sum,
    output logic [31:0] eq
)

endmodule
